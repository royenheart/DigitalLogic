`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 谢皓泽
// 
// Create Date: 2021/10/29 01:44:46
// Design Name: 
// Module Name: ALU32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// 超前进位加法器（32位直接运算）
module G_FullAdder32(
        input wire [31:0]    In1,
        input wire [31:0]    In2,
        input wire           CI,
        input wire           Enable, // Enable Message, high as enable
        output wire [31:0]   Out,
        output wire          CO
    );

    wire [31:0]      OutTmp;
    wire [31:0]      Gi;
    wire [31:0]      Pi;
    wire [31:0]      COi;
    wire [527:0]     CoElement; // The calculate elements of the COi

    // Calculate Gi

    and (Gi[0],In1[0],In2[0]);
    and (Gi[1],In1[1],In2[1]);
    and (Gi[2],In1[2],In2[2]);
    and (Gi[3],In1[3],In2[3]);
    and (Gi[4],In1[4],In2[4]);
    and (Gi[5],In1[5],In2[5]);
    and (Gi[6],In1[6],In2[6]);
    and (Gi[7],In1[7],In2[7]);
    and (Gi[8],In1[8],In2[8]);
    and (Gi[9],In1[9],In2[9]);
    and (Gi[10],In1[10],In2[10]);
    and (Gi[11],In1[11],In2[11]);
    and (Gi[12],In1[12],In2[12]);
    and (Gi[13],In1[13],In2[13]);
    and (Gi[14],In1[14],In2[14]);
    and (Gi[15],In1[15],In2[15]);
    and (Gi[16],In1[16],In2[16]);
    and (Gi[17],In1[17],In2[17]);
    and (Gi[18],In1[18],In2[18]);
    and (Gi[19],In1[19],In2[19]);
    and (Gi[20],In1[20],In2[20]);
    and (Gi[21],In1[21],In2[21]);
    and (Gi[22],In1[22],In2[22]);
    and (Gi[23],In1[23],In2[23]);
    and (Gi[24],In1[24],In2[24]);
    and (Gi[25],In1[25],In2[25]);
    and (Gi[26],In1[26],In2[26]);
    and (Gi[27],In1[27],In2[27]);
    and (Gi[28],In1[28],In2[28]);
    and (Gi[29],In1[29],In2[29]);
    and (Gi[30],In1[30],In2[30]);
    and (Gi[31],In1[31],In2[31]);

    // Calculate Pi

    or (Pi[0],In1[0],In2[0]);
    or (Pi[1],In1[1],In2[1]);
    or (Pi[2],In1[2],In2[2]);
    or (Pi[3],In1[3],In2[3]);
    or (Pi[4],In1[4],In2[4]);
    or (Pi[5],In1[5],In2[5]);
    or (Pi[6],In1[6],In2[6]);
    or (Pi[7],In1[7],In2[7]);
    or (Pi[8],In1[8],In2[8]);
    or (Pi[9],In1[9],In2[9]);
    or (Pi[10],In1[10],In2[10]);
    or (Pi[11],In1[11],In2[11]);
    or (Pi[12],In1[12],In2[12]);
    or (Pi[13],In1[13],In2[13]);
    or (Pi[14],In1[14],In2[14]);
    or (Pi[15],In1[15],In2[15]);
    or (Pi[16],In1[16],In2[16]);
    or (Pi[17],In1[17],In2[17]);
    or (Pi[18],In1[18],In2[18]);
    or (Pi[19],In1[19],In2[19]);
    or (Pi[20],In1[20],In2[20]);
    or (Pi[21],In1[21],In2[21]);
    or (Pi[22],In1[22],In2[22]);
    or (Pi[23],In1[23],In2[23]);
    or (Pi[24],In1[24],In2[24]);
    or (Pi[25],In1[25],In2[25]);
    or (Pi[26],In1[26],In2[26]);
    or (Pi[27],In1[27],In2[27]);
    or (Pi[28],In1[28],In2[28]);
    or (Pi[29],In1[29],In2[29]);
    or (Pi[30],In1[30],In2[30]);
    or (Pi[31],In1[31],In2[31]);

    // Calculate COi's or elements

    and (CoElement[1],Pi[1],Gi[0]);
    and (CoElement[2],CI,Pi[1],Pi[0]);
    and (CoElement[3],Pi[2],Gi[1]);
    and (CoElement[4],Pi[2],Pi[1],Gi[0]);
    and (CoElement[5],CI,Pi[2],Pi[1],Pi[0]);
    and (CoElement[6],Pi[3],Gi[2]);
    and (CoElement[7],Pi[3],Pi[2],Gi[1]);
    and (CoElement[8],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[9],CI,Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[10],Pi[4],Gi[3]);
    and (CoElement[11],Pi[4],Pi[3],Gi[2]);
    and (CoElement[12],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[13],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[14],CI,Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[15],Pi[5],Gi[4]);
    and (CoElement[16],Pi[5],Pi[4],Gi[3]);
    and (CoElement[17],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[18],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[19],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[20],CI,Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[21],Pi[6],Gi[5]);
    and (CoElement[22],Pi[6],Pi[5],Gi[4]);
    and (CoElement[23],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[24],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[25],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[26],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[27],CI,Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[28],Pi[7],Gi[6]);
    and (CoElement[29],Pi[7],Pi[6],Gi[5]);
    and (CoElement[30],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[31],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[32],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[33],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[34],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[35],CI,Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[36],Pi[8],Gi[7]);
    and (CoElement[37],Pi[8],Pi[7],Gi[6]);
    and (CoElement[38],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[39],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[40],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[41],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[42],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[43],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[44],CI,Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[45],Pi[9],Gi[8]);
    and (CoElement[46],Pi[9],Pi[8],Gi[7]);
    and (CoElement[47],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[48],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[49],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[50],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[51],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[52],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[53],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[54],CI,Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[55],Pi[10],Gi[9]);
    and (CoElement[56],Pi[10],Pi[9],Gi[8]);
    and (CoElement[57],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[58],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[59],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[60],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[61],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[62],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[63],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[64],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[65],CI,Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[66],Pi[11],Gi[10]);
    and (CoElement[67],Pi[11],Pi[10],Gi[9]);
    and (CoElement[68],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[69],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[70],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[71],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[72],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[73],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[74],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[75],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[76],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[77],CI,Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[78],Pi[12],Gi[11]);
    and (CoElement[79],Pi[12],Pi[11],Gi[10]);
    and (CoElement[80],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[81],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[82],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[83],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[84],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[85],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[86],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[87],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[88],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[89],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[90],CI,Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[91],Pi[13],Gi[12]);
    and (CoElement[92],Pi[13],Pi[12],Gi[11]);
    and (CoElement[93],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[94],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[95],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[96],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[97],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[98],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[99],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[100],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[101],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[102],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[103],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[104],CI,Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[105],Pi[14],Gi[13]);
    and (CoElement[106],Pi[14],Pi[13],Gi[12]);
    and (CoElement[107],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[108],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[109],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[110],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[111],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[112],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[113],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[114],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[115],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[116],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[117],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[118],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[119],CI,Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[120],Pi[15],Gi[14]);
    and (CoElement[121],Pi[15],Pi[14],Gi[13]);
    and (CoElement[122],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[123],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[124],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[125],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[126],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[127],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[128],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[129],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[130],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[131],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[132],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[133],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[134],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[135],CI,Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[136],Pi[16],Gi[15]);
    and (CoElement[137],Pi[16],Pi[15],Gi[14]);
    and (CoElement[138],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[139],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[140],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[141],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[142],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[143],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[144],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[145],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[146],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[147],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[148],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[149],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[150],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[151],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[152],CI,Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[153],Pi[17],Gi[16]);
    and (CoElement[154],Pi[17],Pi[16],Gi[15]);
    and (CoElement[155],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[156],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[157],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[158],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[159],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[160],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[161],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[162],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[163],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[164],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[165],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[166],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[167],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[168],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[169],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[170],CI,Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[171],Pi[18],Gi[17]);
    and (CoElement[172],Pi[18],Pi[17],Gi[16]);
    and (CoElement[173],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[174],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[175],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[176],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[177],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[178],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[179],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[180],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[181],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[182],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[183],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[184],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[185],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[186],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[187],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[188],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[189],CI,Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[190],Pi[19],Gi[18]);
    and (CoElement[191],Pi[19],Pi[18],Gi[17]);
    and (CoElement[192],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[193],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[194],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[195],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[196],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[197],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[198],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[199],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[200],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[201],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[202],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[203],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[204],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[205],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[206],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[207],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[208],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[209],CI,Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[210],Pi[20],Gi[19]);
    and (CoElement[211],Pi[20],Pi[19],Gi[18]);
    and (CoElement[212],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[213],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[214],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[215],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[216],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[217],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[218],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[219],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[220],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[221],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[222],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[223],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[224],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[225],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[226],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[227],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[228],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[229],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[230],CI,Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[231],Pi[21],Gi[20]);
    and (CoElement[232],Pi[21],Pi[20],Gi[19]);
    and (CoElement[233],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[234],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[235],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[236],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[237],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[238],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[239],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[240],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[241],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[242],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[243],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[244],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[245],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[246],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[247],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[248],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[249],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[250],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[251],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[252],CI,Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[253],Pi[22],Gi[21]);
    and (CoElement[254],Pi[22],Pi[21],Gi[20]);
    and (CoElement[255],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[256],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[257],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[258],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[259],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[260],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[261],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[262],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[263],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[264],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[265],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[266],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[267],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[268],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[269],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[270],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[271],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[272],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[273],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[274],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[275],CI,Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[276],Pi[23],Gi[22]);
    and (CoElement[277],Pi[23],Pi[22],Gi[21]);
    and (CoElement[278],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[279],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[280],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[281],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[282],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[283],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[284],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[285],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[286],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[287],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[288],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[289],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[290],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[291],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[292],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[293],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[294],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[295],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[296],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[297],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[298],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[299],CI,Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[300],Pi[24],Gi[23]);
    and (CoElement[301],Pi[24],Pi[23],Gi[22]);
    and (CoElement[302],Pi[24],Pi[23],Pi[22],Gi[21]);
    and (CoElement[303],Pi[24],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[304],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[305],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[306],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[307],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[308],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[309],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[310],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[311],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[312],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[313],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[314],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[315],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[316],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[317],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[318],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[319],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[320],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[321],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[322],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[323],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[324],CI,Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[325],Pi[25],Gi[24]);
    and (CoElement[326],Pi[25],Pi[24],Gi[23]);
    and (CoElement[327],Pi[25],Pi[24],Pi[23],Gi[22]);
    and (CoElement[328],Pi[25],Pi[24],Pi[23],Pi[22],Gi[21]);
    and (CoElement[329],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[330],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[331],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[332],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[333],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[334],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[335],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[336],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[337],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[338],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[339],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[340],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[341],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[342],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[343],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[344],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[345],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[346],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[347],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[348],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[349],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[350],CI,Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[351],Pi[26],Gi[25]);
    and (CoElement[352],Pi[26],Pi[25],Gi[24]);
    and (CoElement[353],Pi[26],Pi[25],Pi[24],Gi[23]);
    and (CoElement[354],Pi[26],Pi[25],Pi[24],Pi[23],Gi[22]);
    and (CoElement[355],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Gi[21]);
    and (CoElement[356],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[357],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[358],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[359],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[360],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[361],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[362],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[363],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[364],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[365],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[366],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[367],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[368],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[369],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[370],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[371],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[372],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[373],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[374],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[375],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[376],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[377],CI,Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[378],Pi[27],Gi[26]);
    and (CoElement[379],Pi[27],Pi[26],Gi[25]);
    and (CoElement[380],Pi[27],Pi[26],Pi[25],Gi[24]);
    and (CoElement[381],Pi[27],Pi[26],Pi[25],Pi[24],Gi[23]);
    and (CoElement[382],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Gi[22]);
    and (CoElement[383],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Gi[21]);
    and (CoElement[384],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[385],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[386],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[387],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[388],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[389],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[390],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[391],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[392],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[393],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[394],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[395],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[396],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[397],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[398],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[399],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[400],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[401],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[402],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[403],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[404],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[405],CI,Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[406],Pi[28],Gi[27]);
    and (CoElement[407],Pi[28],Pi[27],Gi[26]);
    and (CoElement[408],Pi[28],Pi[27],Pi[26],Gi[25]);
    and (CoElement[409],Pi[28],Pi[27],Pi[26],Pi[25],Gi[24]);
    and (CoElement[410],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Gi[23]);
    and (CoElement[411],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Gi[22]);
    and (CoElement[412],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Gi[21]);
    and (CoElement[413],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[414],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[415],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[416],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[417],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[418],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[419],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[420],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[421],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[422],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[423],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[424],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[425],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[426],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[427],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[428],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[429],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[430],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[431],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[432],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[433],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[434],CI,Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[435],Pi[29],Gi[28]);
    and (CoElement[436],Pi[29],Pi[28],Gi[27]);
    and (CoElement[437],Pi[29],Pi[28],Pi[27],Gi[26]);
    and (CoElement[438],Pi[29],Pi[28],Pi[27],Pi[26],Gi[25]);
    and (CoElement[439],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Gi[24]);
    and (CoElement[440],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Gi[23]);
    and (CoElement[441],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Gi[22]);
    and (CoElement[442],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Gi[21]);
    and (CoElement[443],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[444],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[445],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[446],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[447],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[448],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[449],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[450],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[451],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[452],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[453],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[454],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[455],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[456],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[457],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[458],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[459],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[460],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[461],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[462],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[463],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[464],CI,Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[465],Pi[30],Gi[29]);
    and (CoElement[466],Pi[30],Pi[29],Gi[28]);
    and (CoElement[467],Pi[30],Pi[29],Pi[28],Gi[27]);
    and (CoElement[468],Pi[30],Pi[29],Pi[28],Pi[27],Gi[26]);
    and (CoElement[469],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Gi[25]);
    and (CoElement[470],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Gi[24]);
    and (CoElement[471],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Gi[23]);
    and (CoElement[472],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Gi[22]);
    and (CoElement[473],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Gi[21]);
    and (CoElement[474],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[475],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[476],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[477],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[478],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[479],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[480],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[481],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[482],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[483],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[484],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[485],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[486],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[487],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[488],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[489],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[490],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[491],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[492],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[493],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[494],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[495],CI,Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);
    and (CoElement[496],Pi[31],Gi[30]);
    and (CoElement[497],Pi[31],Pi[30],Gi[29]);
    and (CoElement[498],Pi[31],Pi[30],Pi[29],Gi[28]);
    and (CoElement[499],Pi[31],Pi[30],Pi[29],Pi[28],Gi[27]);
    and (CoElement[500],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Gi[26]);
    and (CoElement[501],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Gi[25]);
    and (CoElement[502],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Gi[24]);
    and (CoElement[503],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Gi[23]);
    and (CoElement[504],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Gi[22]);
    and (CoElement[505],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Gi[21]);
    and (CoElement[506],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Gi[20]);
    and (CoElement[507],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Gi[19]);
    and (CoElement[508],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Gi[18]);
    and (CoElement[509],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Gi[17]);
    and (CoElement[510],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Gi[16]);
    and (CoElement[511],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Gi[15]);
    and (CoElement[512],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Gi[14]);
    and (CoElement[513],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Gi[13]);
    and (CoElement[514],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Gi[12]);
    and (CoElement[515],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Gi[11]);
    and (CoElement[516],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Gi[10]);
    and (CoElement[517],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Gi[9]);
    and (CoElement[518],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Gi[8]);
    and (CoElement[519],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Gi[7]);
    and (CoElement[520],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Gi[6]);
    and (CoElement[521],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Gi[5]);
    and (CoElement[522],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Gi[4]);
    and (CoElement[523],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Gi[3]);
    and (CoElement[524],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Gi[2]);
    and (CoElement[525],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Gi[1]);
    and (CoElement[526],Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Gi[0]);
    and (CoElement[527],CI,Pi[31],Pi[30],Pi[29],Pi[28],Pi[27],Pi[26],Pi[25],Pi[24],Pi[23],Pi[22],Pi[21],Pi[20],Pi[19],Pi[18],Pi[17],Pi[16],Pi[15],Pi[14],Pi[13],Pi[12],Pi[11],Pi[10],Pi[9],Pi[8],Pi[7],Pi[6],Pi[5],Pi[4],Pi[3],Pi[2],Pi[1],Pi[0]);


    // Calculate COi

    or (COi[0],Gi[0],CoElement[0]);
    or (COi[1],Gi[1],CoElement[2],CoElement[1]);
    or (COi[2],Gi[2],CoElement[5],CoElement[4],CoElement[3]);
    or (COi[3],Gi[3],CoElement[9],CoElement[8],CoElement[7],CoElement[6]);
    or (COi[4],Gi[4],CoElement[14],CoElement[13],CoElement[12],CoElement[11],CoElement[10]);
    or (COi[5],Gi[5],CoElement[20],CoElement[19],CoElement[18],CoElement[17],CoElement[16],CoElement[15]);
    or (COi[6],Gi[6],CoElement[27],CoElement[26],CoElement[25],CoElement[24],CoElement[23],CoElement[22],CoElement[21]);
    or (COi[7],Gi[7],CoElement[35],CoElement[34],CoElement[33],CoElement[32],CoElement[31],CoElement[30],CoElement[29],CoElement[28]);
    or (COi[8],Gi[8],CoElement[44],CoElement[43],CoElement[42],CoElement[41],CoElement[40],CoElement[39],CoElement[38],CoElement[37],CoElement[36]);
    or (COi[9],Gi[9],CoElement[54],CoElement[53],CoElement[52],CoElement[51],CoElement[50],CoElement[49],CoElement[48],CoElement[47],CoElement[46],CoElement[45]);
    or (COi[10],Gi[10],CoElement[65],CoElement[64],CoElement[63],CoElement[62],CoElement[61],CoElement[60],CoElement[59],CoElement[58],CoElement[57],CoElement[56],CoElement[55]);
    or (COi[11],Gi[11],CoElement[77],CoElement[76],CoElement[75],CoElement[74],CoElement[73],CoElement[72],CoElement[71],CoElement[70],CoElement[69],CoElement[68],CoElement[67],CoElement[66]);
    or (COi[12],Gi[12],CoElement[90],CoElement[89],CoElement[88],CoElement[87],CoElement[86],CoElement[85],CoElement[84],CoElement[83],CoElement[82],CoElement[81],CoElement[80],CoElement[79],CoElement[78]);
    or (COi[13],Gi[13],CoElement[104],CoElement[103],CoElement[102],CoElement[101],CoElement[100],CoElement[99],CoElement[98],CoElement[97],CoElement[96],CoElement[95],CoElement[94],CoElement[93],CoElement[92],CoElement[91]);
    or (COi[14],Gi[14],CoElement[119],CoElement[118],CoElement[117],CoElement[116],CoElement[115],CoElement[114],CoElement[113],CoElement[112],CoElement[111],CoElement[110],CoElement[109],CoElement[108],CoElement[107],CoElement[106],CoElement[105]);
    or (COi[15],Gi[15],CoElement[135],CoElement[134],CoElement[133],CoElement[132],CoElement[131],CoElement[130],CoElement[129],CoElement[128],CoElement[127],CoElement[126],CoElement[125],CoElement[124],CoElement[123],CoElement[122],CoElement[121],CoElement[120]);
    or (COi[16],Gi[16],CoElement[152],CoElement[151],CoElement[150],CoElement[149],CoElement[148],CoElement[147],CoElement[146],CoElement[145],CoElement[144],CoElement[143],CoElement[142],CoElement[141],CoElement[140],CoElement[139],CoElement[138],CoElement[137],CoElement[136]);
    or (COi[17],Gi[17],CoElement[170],CoElement[169],CoElement[168],CoElement[167],CoElement[166],CoElement[165],CoElement[164],CoElement[163],CoElement[162],CoElement[161],CoElement[160],CoElement[159],CoElement[158],CoElement[157],CoElement[156],CoElement[155],CoElement[154],CoElement[153]);
    or (COi[18],Gi[18],CoElement[189],CoElement[188],CoElement[187],CoElement[186],CoElement[185],CoElement[184],CoElement[183],CoElement[182],CoElement[181],CoElement[180],CoElement[179],CoElement[178],CoElement[177],CoElement[176],CoElement[175],CoElement[174],CoElement[173],CoElement[172],CoElement[171]);
    or (COi[19],Gi[19],CoElement[209],CoElement[208],CoElement[207],CoElement[206],CoElement[205],CoElement[204],CoElement[203],CoElement[202],CoElement[201],CoElement[200],CoElement[199],CoElement[198],CoElement[197],CoElement[196],CoElement[195],CoElement[194],CoElement[193],CoElement[192],CoElement[191],CoElement[190]);
    or (COi[20],Gi[20],CoElement[230],CoElement[229],CoElement[228],CoElement[227],CoElement[226],CoElement[225],CoElement[224],CoElement[223],CoElement[222],CoElement[221],CoElement[220],CoElement[219],CoElement[218],CoElement[217],CoElement[216],CoElement[215],CoElement[214],CoElement[213],CoElement[212],CoElement[211],CoElement[210]);
    or (COi[21],Gi[21],CoElement[252],CoElement[251],CoElement[250],CoElement[249],CoElement[248],CoElement[247],CoElement[246],CoElement[245],CoElement[244],CoElement[243],CoElement[242],CoElement[241],CoElement[240],CoElement[239],CoElement[238],CoElement[237],CoElement[236],CoElement[235],CoElement[234],CoElement[233],CoElement[232],CoElement[231]);
    or (COi[22],Gi[22],CoElement[275],CoElement[274],CoElement[273],CoElement[272],CoElement[271],CoElement[270],CoElement[269],CoElement[268],CoElement[267],CoElement[266],CoElement[265],CoElement[264],CoElement[263],CoElement[262],CoElement[261],CoElement[260],CoElement[259],CoElement[258],CoElement[257],CoElement[256],CoElement[255],CoElement[254],CoElement[253]);
    or (COi[23],Gi[23],CoElement[299],CoElement[298],CoElement[297],CoElement[296],CoElement[295],CoElement[294],CoElement[293],CoElement[292],CoElement[291],CoElement[290],CoElement[289],CoElement[288],CoElement[287],CoElement[286],CoElement[285],CoElement[284],CoElement[283],CoElement[282],CoElement[281],CoElement[280],CoElement[279],CoElement[278],CoElement[277],CoElement[276]);
    or (COi[24],Gi[24],CoElement[324],CoElement[323],CoElement[322],CoElement[321],CoElement[320],CoElement[319],CoElement[318],CoElement[317],CoElement[316],CoElement[315],CoElement[314],CoElement[313],CoElement[312],CoElement[311],CoElement[310],CoElement[309],CoElement[308],CoElement[307],CoElement[306],CoElement[305],CoElement[304],CoElement[303],CoElement[302],CoElement[301],CoElement[300]);
    or (COi[25],Gi[25],CoElement[350],CoElement[349],CoElement[348],CoElement[347],CoElement[346],CoElement[345],CoElement[344],CoElement[343],CoElement[342],CoElement[341],CoElement[340],CoElement[339],CoElement[338],CoElement[337],CoElement[336],CoElement[335],CoElement[334],CoElement[333],CoElement[332],CoElement[331],CoElement[330],CoElement[329],CoElement[328],CoElement[327],CoElement[326],CoElement[325]);
    or (COi[26],Gi[26],CoElement[377],CoElement[376],CoElement[375],CoElement[374],CoElement[373],CoElement[372],CoElement[371],CoElement[370],CoElement[369],CoElement[368],CoElement[367],CoElement[366],CoElement[365],CoElement[364],CoElement[363],CoElement[362],CoElement[361],CoElement[360],CoElement[359],CoElement[358],CoElement[357],CoElement[356],CoElement[355],CoElement[354],CoElement[353],CoElement[352],CoElement[351]);
    or (COi[27],Gi[27],CoElement[405],CoElement[404],CoElement[403],CoElement[402],CoElement[401],CoElement[400],CoElement[399],CoElement[398],CoElement[397],CoElement[396],CoElement[395],CoElement[394],CoElement[393],CoElement[392],CoElement[391],CoElement[390],CoElement[389],CoElement[388],CoElement[387],CoElement[386],CoElement[385],CoElement[384],CoElement[383],CoElement[382],CoElement[381],CoElement[380],CoElement[379],CoElement[378]);
    or (COi[28],Gi[28],CoElement[434],CoElement[433],CoElement[432],CoElement[431],CoElement[430],CoElement[429],CoElement[428],CoElement[427],CoElement[426],CoElement[425],CoElement[424],CoElement[423],CoElement[422],CoElement[421],CoElement[420],CoElement[419],CoElement[418],CoElement[417],CoElement[416],CoElement[415],CoElement[414],CoElement[413],CoElement[412],CoElement[411],CoElement[410],CoElement[409],CoElement[408],CoElement[407],CoElement[406]);
    or (COi[29],Gi[29],CoElement[464],CoElement[463],CoElement[462],CoElement[461],CoElement[460],CoElement[459],CoElement[458],CoElement[457],CoElement[456],CoElement[455],CoElement[454],CoElement[453],CoElement[452],CoElement[451],CoElement[450],CoElement[449],CoElement[448],CoElement[447],CoElement[446],CoElement[445],CoElement[444],CoElement[443],CoElement[442],CoElement[441],CoElement[440],CoElement[439],CoElement[438],CoElement[437],CoElement[436],CoElement[435]);
    or (COi[30],Gi[30],CoElement[495],CoElement[494],CoElement[493],CoElement[492],CoElement[491],CoElement[490],CoElement[489],CoElement[488],CoElement[487],CoElement[486],CoElement[485],CoElement[484],CoElement[483],CoElement[482],CoElement[481],CoElement[480],CoElement[479],CoElement[478],CoElement[477],CoElement[476],CoElement[475],CoElement[474],CoElement[473],CoElement[472],CoElement[471],CoElement[470],CoElement[469],CoElement[468],CoElement[467],CoElement[466],CoElement[465]);
    or (COi[31],Gi[31],CoElement[527],CoElement[526],CoElement[525],CoElement[524],CoElement[523],CoElement[522],CoElement[521],CoElement[520],CoElement[519],CoElement[518],CoElement[517],CoElement[516],CoElement[515],CoElement[514],CoElement[513],CoElement[512],CoElement[511],CoElement[510],CoElement[509],CoElement[508],CoElement[507],CoElement[506],CoElement[505],CoElement[504],CoElement[503],CoElement[502],CoElement[501],CoElement[500],CoElement[499],CoElement[498],CoElement[497],CoElement[496]);
    buf     (CO,COi[31]);

    // Calculate Out 

    xor (Out[0],In1[0],In2[0],CI);
    xor (Out[1],In1[1],In2[1],COi[0]);    
    xor (Out[2],In1[2],In2[2],COi[1]);    
    xor (Out[3],In1[3],In2[3],COi[2]);    
    xor (Out[4],In1[4],In2[4],COi[3]);    
    xor (Out[5],In1[5],In2[5],COi[4]);    
    xor (Out[6],In1[6],In2[6],COi[5]);    
    xor (Out[7],In1[7],In2[7],COi[6]);    
    xor (Out[8],In1[8],In2[8],COi[7]);    
    xor (Out[9],In1[9],In2[9],COi[8]);    
    xor (Out[10],In1[10],In2[10],COi[9]); 
    xor (Out[11],In1[11],In2[11],COi[10]);
    xor (Out[12],In1[12],In2[12],COi[11]);
    xor (Out[13],In1[13],In2[13],COi[12]);
    xor (Out[14],In1[14],In2[14],COi[13]);
    xor (Out[15],In1[15],In2[15],COi[14]);
    xor (Out[16],In1[16],In2[16],COi[15]);
    xor (Out[17],In1[17],In2[17],COi[16]);
    xor (Out[18],In1[18],In2[18],COi[17]);
    xor (Out[19],In1[19],In2[19],COi[18]);
    xor (Out[20],In1[20],In2[20],COi[19]);
    xor (Out[21],In1[21],In2[21],COi[20]);
    xor (Out[22],In1[22],In2[22],COi[21]);
    xor (Out[23],In1[23],In2[23],COi[22]);
    xor (Out[24],In1[24],In2[24],COi[23]);
    xor (Out[25],In1[25],In2[25],COi[24]);
    xor (Out[26],In1[26],In2[26],COi[25]);
    xor (Out[27],In1[27],In2[27],COi[26]);
    xor (Out[28],In1[28],In2[28],COi[27]);
    xor (Out[29],In1[29],In2[29],COi[28]);
    xor (Out[30],In1[30],In2[30],COi[29]);
    xor (Out[31],In1[31],In2[31],COi[30]);

    // And Enable Message to Out

    and     (Out[0],OutTmp[0],Enable);
    and     (Out[1],OutTmp[1],Enable);
    and     (Out[2],OutTmp[2],Enable);
    and     (Out[3],OutTmp[3],Enable);
    and     (Out[4],OutTmp[4],Enable);
    and     (Out[5],OutTmp[5],Enable);
    and     (Out[6],OutTmp[6],Enable);
    and     (Out[7],OutTmp[7],Enable);
    and     (Out[8],OutTmp[8],Enable);
    and     (Out[9],OutTmp[9],Enable);
    and     (Out[10],OutTmp[10],Enable);
    and     (Out[11],OutTmp[11],Enable);
    and     (Out[12],OutTmp[12],Enable);
    and     (Out[13],OutTmp[13],Enable);
    and     (Out[14],OutTmp[14],Enable);
    and     (Out[15],OutTmp[15],Enable);
    and     (Out[16],OutTmp[16],Enable);
    and     (Out[17],OutTmp[17],Enable);
    and     (Out[18],OutTmp[18],Enable);
    and     (Out[19],OutTmp[19],Enable);
    and     (Out[20],OutTmp[20],Enable);
    and     (Out[21],OutTmp[21],Enable);
    and     (Out[22],OutTmp[22],Enable);
    and     (Out[23],OutTmp[23],Enable);
    and     (Out[24],OutTmp[24],Enable);
    and     (Out[25],OutTmp[25],Enable);
    and     (Out[26],OutTmp[26],Enable);
    and     (Out[27],OutTmp[27],Enable);
    and     (Out[28],OutTmp[28],Enable);
    and     (Out[29],OutTmp[29],Enable);
    and     (Out[30],OutTmp[30],Enable);
    and     (Out[31],OutTmp[31],Enable);

endmodule