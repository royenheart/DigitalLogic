`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 
// Design Name: 
// Module Name: FFT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 使用FFT快速傅里叶变换+蝴蝶操作对2个1024位大数进行乘法运算
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Addi    tional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module FFT (
    input wire [1023:0] In1,
    input wire [1023:0] In2
);
    
endmodule