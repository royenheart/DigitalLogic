`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 谢皓泽
// 
// Create Date: 2021/10/28 15:52:59
// Design Name: 
// Module Name: And32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// RTL级32位高、低位截断
module Truncated (
        input wire [31:0]  In1,
        input wire [31:0]  In2,
        output wire [31:0] Out
    );

    reg [31:0] tmp;
    reg  i;

    assign  Out = tmp;

    always @(*) 
    begin
        case (In2[31])
            1'b1: 
            begin
                tmp = ( In1 << (32-In2[4:0]) ) >> (32-In2[4:0]);
            end
            1'b0: 
            begin
                tmp = ( In1 >> (32-In2[4:0]) );
            end
            default: tmp = 0;
        endcase    
    end

endmodule
